** Profile: "Z-Measurement-Setup-Profile1"  [ c:\dev\tauv-hardware\tauv-acoustics-v2\simulation\transducer-characterization\transducer-characterization-pspicefiles\z-measurement-setup\profile1.sim ] 

** Creating circuit file "Profile1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Gleb Ryabtsev\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1k 10Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Z-Measurement-Setup.net" 


.END
